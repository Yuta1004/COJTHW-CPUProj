module cpu_core_controller_v1_0 #
    (
        parameter integer C_S_AXI_DATA_WIDTH    = 32,
        parameter integer C_S_AXI_ADDR_WIDTH    = 16
    )
    (
        // CORE�Ƃ̐ڑ��|�[�g
        input wire          CCLK,
        output wire         CRST,
        input wire [31:0]   REG00,
        input wire [31:0]   REG01,
        input wire [31:0]   REG02,
        input wire [31:0]   REG03,
        input wire [31:0]   REG04,
        input wire [31:0]   REG05,
        input wire [31:0]   REG06,
        input wire [31:0]   REG07,
        input wire [31:0]   REG08,
        input wire [31:0]   REG09,
        input wire [31:0]   REG10,
        input wire [31:0]   REG11,
        input wire [31:0]   REG12,
        input wire [31:0]   REG13,
        input wire [31:0]   REG14,
        input wire [31:0]   REG15,
        input wire [31:0]   REG16,
        input wire [31:0]   REG17,
        input wire [31:0]   REG18,
        input wire [31:0]   REG19,
        input wire [31:0]   REG20,
        input wire [31:0]   REG21,
        input wire [31:0]   REG22,
        input wire [31:0]   REG23,
        input wire [31:0]   REG24,
        input wire [31:0]   REG25,
        input wire [31:0]   REG26,
        input wire [31:0]   REG27,
        input wire [31:0]   REG28,
        input wire [31:0]   REG29,
        input wire [31:0]   REG30,
        input wire [31:0]   REG31,
        input wire [31:0]   REGPC,

        input wire  s_axi_aclk,
        input wire  s_axi_aresetn,
        input wire [C_S_AXI_ADDR_WIDTH-1 : 0] s_axi_awaddr,
        input wire [2 : 0] s_axi_awprot,
        input wire  s_axi_awvalid,
        output wire  s_axi_awready,
        input wire [C_S_AXI_DATA_WIDTH-1 : 0] s_axi_wdata,
        input wire [(C_S_AXI_DATA_WIDTH/8)-1 : 0] s_axi_wstrb,
        input wire  s_axi_wvalid,
        output wire  s_axi_wready,
        output wire [1 : 0] s_axi_bresp,
        output wire  s_axi_bvalid,
        input wire  s_axi_bready,
        input wire [C_S_AXI_ADDR_WIDTH-1 : 0] s_axi_araddr,
        input wire [2 : 0] s_axi_arprot,
        input wire  s_axi_arvalid,
        output wire  s_axi_arready,
        output wire [C_S_AXI_DATA_WIDTH-1 : 0] s_axi_rdata,
        output wire [1 : 0] s_axi_rresp,
        output wire  s_axi_rvalid,
        input wire  s_axi_rready
    );

    cpu_core_controller_v1_0_S_AXI # (
        .C_S_AXI_DATA_WIDTH(C_S_AXI_DATA_WIDTH),
        .C_S_AXI_ADDR_WIDTH(C_S_AXI_ADDR_WIDTH)
    ) cpu_core_controller_v1_0_S_AXI_inst (
        .CCLK(CCLK),
        .CRST(CRST),
        .REG00(REG00),
        .REG01(REG01),
        .REG02(REG02),
        .REG03(REG03),
        .REG04(REG04),
        .REG05(REG05),
        .REG06(REG06),
        .REG07(REG07),
        .REG08(REG08),
        .REG09(REG09),
        .REG10(REG10),
        .REG11(REG11),
        .REG12(REG12),
        .REG13(REG13),
        .REG14(REG14),
        .REG15(REG15),
        .REG16(REG16),
        .REG17(REG17),
        .REG18(REG18),
        .REG19(REG19),
        .REG20(REG20),
        .REG21(REG21),
        .REG22(REG22),
        .REG23(REG23),
        .REG24(REG24),
        .REG25(REG25),
        .REG26(REG26),
        .REG27(REG27),
        .REG28(REG28),
        .REG29(REG229),
        .REG30(REG30),
        .REG31(REG31),
        .REGPC(REGPC),
        .S_AXI_ACLK(s_axi_aclk),
        .S_AXI_ARESETN(s_axi_aresetn),
        .S_AXI_AWADDR(s_axi_awaddr),
        .S_AXI_AWPROT(s_axi_awprot),
        .S_AXI_AWVALID(s_axi_awvalid),
        .S_AXI_AWREADY(s_axi_awready),
        .S_AXI_WDATA(s_axi_wdata),
        .S_AXI_WSTRB(s_axi_wstrb),
        .S_AXI_WVALID(s_axi_wvalid),
        .S_AXI_WREADY(s_axi_wready),
        .S_AXI_BRESP(s_axi_bresp),
        .S_AXI_BVALID(s_axi_bvalid),
        .S_AXI_BREADY(s_axi_bready),
        .S_AXI_ARADDR(s_axi_araddr),
        .S_AXI_ARPROT(s_axi_arprot),
        .S_AXI_ARVALID(s_axi_arvalid),
        .S_AXI_ARREADY(s_axi_arready),
        .S_AXI_RDATA(s_axi_rdata),
        .S_AXI_RRESP(s_axi_rresp),
        .S_AXI_RVALID(s_axi_rvalid),
        .S_AXI_RREADY(s_axi_rready)
    );

endmodule
